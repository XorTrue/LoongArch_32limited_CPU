`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/07/23 20:15:46
// Design Name: 
// Module Name: ID_EX0
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ID_EX0(
    input clk, rst,

    input ID_EX0_stall_from_DCache,
    input ID_EX0_flush_from_EX_Branch


    );
endmodule
